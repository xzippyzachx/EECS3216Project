module EECS3216Project ();
	
	
endmodule